module iopoller


fn test_1() {
    
}
