module corona

fn test_compile() {

}

